module top(
    input [7:0] in,
    input clk,
    output [7:0] out
    );
    
    //Add code here

    
endmodule
